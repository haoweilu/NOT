module NOT(
    input a,
    output b
);

    assign b = ~a;

endmodule